constant rom : integer_array := (0,
0,
0,
0,
0,
1,
1,
1,
1,
0,
-1,
-4,
-7,
-10,
-14,
-16,
-17,
-15,
-10,
0,
15,
35,
59,
87,
116,
143,
168,
188,
201,
205,
201,
188,
168,
143,
116,
87,
59,
35,
15,
0,
-10,
-15,
-17,
-16,
-14,
-10,
-7,
-4,
-1,
0,
1,
1,
1,
1,
0,
0,
0,
0,
0
);