constant rom : integer_array := (0,
0,
1,
1,
1,
0,
-1,
-3,
-4,
-1,
2,
6,
7,
4,
-3,
-9,
-10,
-6,
2,
8,
9,
5,
0,
-2,
0,
3,
1,
-9,
-19,
-21,
-6,
22,
48,
51,
21,
-33,
-80,
-89,
-44,
35,
107,
126,
74,
-27,
-122,
-154,
-101,
10,
119,
2212,
119,
10,
-101,
-153,
-120,
-27,
73,
124,
105,
34,
-44,
-86,
-78,
-32,
20,
49,
46,
21,
-6,
-20,
-18,
-8,
0,
3,
0,
-2,
0,
5,
8,
7,
2,
-5,
-9,
-8,
-3,
3,
6,
6,
2,
-1,
-3,
-3,
-1,
0,
1,
1,
1,
0,
0
);