constant rom : integer_array := (0,
0,
0,
0,
0,
-1,
-1,
-1,
-1,
-1,
-2,
-2,
-2,
-2,
-2,
-2,
6132,
-2,
-2,
-2,
-2,
-2,
-1,
-1,
-1,
-1,
-1,
0,
0,
0,
0,
0,
0
);